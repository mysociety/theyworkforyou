2004-01-19
Leader|Ian Paisley
Deputy Leader|Peter Robinson
Whip|Nigel Dodds
Whip|Gergory Campbell
Whip|Jeffrey Donaldson
Whip|Iris Robinson
2004-12-13
Leader|Ian Paisley
Deputy Leader|Peter Robinson
Whip|Nigel Dodds
Whip|Gergory Campbell
Whip|Jeffrey Donaldson
Whip|Andrew Hunter
Whip|Iris Robinson
2006-04-28
Leader; Foreign & Commonwealth Affairs; Europe|Rt Hon Ian Paisley MP
Deputy Leader; Home Affairs; Constitutional Affairs|Peter Robinson MP
Treasury; Work and Pensions; Shadow Leader of the House|Nigel Dodds MP
Defence; Culture, Media & Sport|Gregory Campbell MP
Transport, International Development|Jeffrey Donaldson MP
Environment, Food & Rural Affairs|Rev Dr William McCrea MP
Health, Youth & Women|Iris Robinson MP
Trade and Industry|David Simpson MP
Education and Skills; Housing (ODPM)|Sammy Wilson MP
2006-08-02
Leader; Foreign & Commonwealth Affairs; Europe|Rt Hon Ian Paisley MP
Deputy Leader; Home Affairs; Constitutional Affairs|Peter Robinson MP
Treasury; Work and Pensions; Shadow Leader of the House|Nigel Dodds MP
Defence; Culture, Media & Sport|Gregory Campbell MP
Transport, International Development|Jeffrey Donaldson MP
Environment, Food & Rural Affairs|Rev Dr William McCrea MP
Health, Youth & Women|Iris Robinson MP
Trade and Industry|David Simpson MP
Education and Skills; Housing (DCLG)|Sammy Wilson MP
2007-05-10
Leader; Foreign & Commonwealth Affairs; Europe|Rt Hon Ian Paisley MP
Deputy Leader; Home Affairs; Constitutional Affairs|Rt Hon Peter Robinson MP
Treasury; Work and Pensions; Shadow Leader of the House|Nigel Dodds MP
Defence; Culture, Media & Sport|Gregory Campbell MP
Transport, International Development|Rt Hon Jeffrey Donaldson MP
Environment, Food & Rural Affairs|Rev Dr William McCrea MP
Health, Youth & Women|Iris Robinson MP
Trade and Industry|David Simpson MP
Education and Skills; Housing (DCLG)|Sammy Wilson MP
2007-07-27
Leader; Foreign & Commonwealth Affairs; Europe|Rt Hon Ian Paisley MP
Deputy Leader; Home Affairs; Constitutional Affairs|Rt Hon Peter Robinson MP
Treasury; Work and Pensions; Shadow Leader of the House|Nigel Dodds MP
Defence; Culture, Media & Sport|Gregory Campbell MP
Transport, International Development|Rt Hon Jeffrey Donaldson MP
Environment, Food & Rural Affairs|Rev Dr William McCrea MP
Health  & Women|Iris Robinson MP
Trade and Industry; Young People|David Simpson MP
Children, Schools and Families; Communities and Local Government|Sammy Wilson MP
